.title KiCad schematic
44B_P10 1 2 3 4 5 3 0 6 3 7 8 3 9 10 7402
33B_P10 3 11 12 13 14 15 0 16 17 10 74HC04
22E_P10 18 19 20 21 22 0 3 23 20 19 18 10 74LS13
22B_P10 24 25 26 6 27 8 0 28 29 30 31 32 33 10 74HC04
22A_P10 34 2 35 36 37 35 0 38 39 40 38 5 41 10 74HC04
11B_P10 42 43 44 45 46 44 0 23 47 21 23 48 43 10 74HC04
11A_P10 49 20 50 19 51 50 0 52 53 18 52 54 20 10 74HC04
44C_P10 55 54 56 57 56 20 0 58 20 59 54 58 60 10 7402
33A_P10 61 62 58 63 56 64 0 65 22 66 67 68 69 10 74HC04
44D_P10 52 21 61 50 52 56 0 58 52 19 10 7400
55C_P10 70 21 67 71 67 23 0 69 23 72 21 69 73 10 7402
11C_P10 18 19 18 50 54 69 0 74 36 40 48 67 54 10 74LS10
55B_P10 75 44 22 76 43 22 0 35 22 77 38 22 78 10 7402
55A_P10 79 80 14 81 82 14 0 83 14 84 85 14 86 10 7402
33C_P10 87 74 14 0 10 7402
44A_P10 88 12 21 89 14 90 0 91 14 92 93 14 94 10 7402
33D_P10 43 38 43 38 36 93 0 91 35 40 43 90 35 10 74LS10
11E_P10 43 40 0 80 36 10 74LS10
22D_P10 48 38 48 38 36 85 0 12 20 50 18 82 35 10 74LS10
11D_P10 13 21 13 21 44 17 0 83 35 40 48 14 45 10 74LS10
22C_P10 2 5 8 6 25 28 0 95 30 32 10 74LS30
CCONECTOR_P10 10 53 51 49 47 46 42 39 37 95 96 97 98 99 100 63 64 68 66 62 65 87 55 57 88 89 1 4 75 76 79 81 70 71 101 102 34 41 27 26 24 29 31 33 52 103 104 105 106 107 11 15 16 13 108 109 110 60 59 94 92 9 7 78 77 86 84 73 72 0 CONN_35X2
.end
